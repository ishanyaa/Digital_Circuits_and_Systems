module or3 (output Y, input A, B, C);

  // Structural description using built-in OR gate
  or (Y, A, B, C);

endmodule
