//Problem 1 A-1

module and3 (output Y, input A, B, C);

and(Y,A,B,);

endmodule